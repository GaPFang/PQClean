`timescale 1ns/1ps

module ntt_tb;

  // Parameters
  localparam [31:0] KYBER_Q = 3329;

  // Clock / reset / control
  logic clk;
  logic rst_n;
  logic ready;
  logic valid;
  logic tmp_valid;
  logic [31:0] i_addr;
  logic [31:0] i_Kyber_ntt_config, i_Kyber_intt_config, i_Dilithium_ntt_config, i_Dilithium_intt_config;
  logic signed [31:0] tmp_data;

  // Input / output arrays (SystemVerilog unpacked arrays)
  logic signed [31:0] i_data;
  logic signed [31:0] o_data;
  logic signed [31:0] r_out [0:255];

  // Instantiate DUT (adjust instance name / port names if your module differs)
  ntt dut_ntt (
    .ntt_clk_i   (clk),
    .ntt_rst_ni  (rst_n),

    .ntt_req_i   (),
    .ntt_we_i    (ready | i_addr[2]),
    .ntt_be_i    (),
    .ntt_addr_i  (i_addr),
    .ntt_wdata_i (i_addr[2] ? i_Dilithium_ntt_config : i_data),
    .ntt_rvalid_o(tmp_valid),
    .ntt_rdata_o (tmp_data),
    .ntt_err_o   (),
    .ntt_intr_o  ()
  );

  ntt dut_intt (
    .ntt_clk_i   (clk),
    .ntt_rst_ni  (rst_n),

    .ntt_req_i   (),
    .ntt_we_i    (tmp_valid | i_addr[2]),
    .ntt_be_i    (),
    .ntt_addr_i  (i_addr),
    .ntt_wdata_i (i_addr[2] ? i_Dilithium_intt_config : tmp_data),
    .ntt_rvalid_o(valid),
    .ntt_rdata_o (o_data),
    .ntt_err_o   (),
    .ntt_intr_o  ()
  );

  integer cycles;

  // Clock generation: 10 ns period
  initial begin
    clk = 0;
    forever #5 clk = ~clk;
  end

  initial begin
    while (1) begin
      @(posedge clk);
      cycles = cycles + 1;
    end
  end

  // Test scenario
  logic [31:0] i;
  initial begin
    $fsdbDumpfile("ntt_tb.fsdb");
    $fsdbDumpvars;
    $fsdbDumpMDA;
    // $dumpfile("ntt_tb.vcd");
    // $dumpvars(0, ntt_tb);

    // Reset
    rst_n = 0;
    ready = 0;
    repeat (4) @(posedge clk);
    rst_n = 1;
    i_data = 0;
    cycles = 0;
    @(posedge clk);
    ready = 1;
    i_addr = 3'b100;
    i_Kyber_ntt_config = 2'b00;
    i_Kyber_intt_config = 2'b01;
    i_Dilithium_ntt_config = 2'b10;
    i_Dilithium_intt_config = 2'b11;
    @(posedge clk);
    i_addr = 0;
    // Step 1: Prepare input like C code: r[i] = i % KYBER_Q
    for (i = 0; i < 256; i = i + 1) begin
      i_data = (i % KYBER_Q); // fits in 16-bit signed
      @(posedge clk);
    end
    ready = 0;
    $display("Input finish: %d cycles", cycles);

    // give one clock to allow o_data to be stable if needed
    @(posedge clk);

    i = 0;
    while (i < 256) begin
      @(negedge clk);
      if (valid) begin
        if (i == 0) begin
          $display("Computation finish: %d cycles", cycles);
        end
        r_out[i] = o_data;
        i = i + 1;
      end
    end

    $display("Output finish: %d cycles", cycles);

    // Step 3: print results, 16 per line like C code
    $display("NTT result:");
    for (i = 0; i < 256; i = i + 1) begin
      // sign-printed decimal with width 6 to mimic printf("%6d ")
      $write("%5d ", $signed(r_out[i]));
      if (((i + 1) % 16) == 0) $write("\n");
    end
    $write("\n");

    // finish
    $display("Test finished.");
    #10;
    $finish;
  end

endmodule
